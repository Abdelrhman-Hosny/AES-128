module AESFull(input a,b, output c);
assign c = a & b;
endmodule