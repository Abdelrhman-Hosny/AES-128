module InvSBox(input clk,input [7:0] input_byte, output reg[7:0] output_byte);
always @(posedge clk) begin
case(input_byte)
8'h63: output_byte = 8'h00;
8'h7c: output_byte = 8'h01;
8'h77: output_byte = 8'h02;
8'h7b: output_byte = 8'h03;
8'hf2: output_byte = 8'h04;
8'h6b: output_byte = 8'h05;
8'h6f: output_byte = 8'h06;
8'hc5: output_byte = 8'h07;
8'h30: output_byte = 8'h08;
8'h01: output_byte = 8'h09;
8'h67: output_byte = 8'h0A;
8'h2b: output_byte = 8'h0B;
8'hfe: output_byte = 8'h0C;
8'hd7: output_byte = 8'h0D;
8'hab: output_byte = 8'h0E;
8'h76: output_byte = 8'h0F;
8'hca: output_byte = 8'h10;
8'h82: output_byte = 8'h11;
8'hc9: output_byte = 8'h12;
8'h7d: output_byte = 8'h13;
8'hfa: output_byte = 8'h14;
8'h59: output_byte = 8'h15;
8'h47: output_byte = 8'h16;
8'hf0: output_byte = 8'h17;
8'had: output_byte = 8'h18;
8'hd4: output_byte = 8'h19;
8'ha2: output_byte = 8'h1A;
8'haf: output_byte = 8'h1B;
8'h9c: output_byte = 8'h1C;
8'ha4: output_byte = 8'h1D;
8'h72: output_byte = 8'h1E;
8'hc0: output_byte = 8'h1F;
8'hb7: output_byte = 8'h20;
8'hfd: output_byte = 8'h21;
8'h93: output_byte = 8'h22;
8'h26: output_byte = 8'h23;
8'h36: output_byte = 8'h24;
8'h3f: output_byte = 8'h25;
8'hf7: output_byte = 8'h26;
8'hcc: output_byte = 8'h27;
8'h34: output_byte = 8'h28;
8'ha5: output_byte = 8'h29;
8'he5: output_byte = 8'h2A;
8'hf1: output_byte = 8'h2B;
8'h71: output_byte = 8'h2C;
8'hd8: output_byte = 8'h2D;
8'h31: output_byte = 8'h2E;
8'h15: output_byte = 8'h2F;
8'h04: output_byte = 8'h30;
8'hc7: output_byte = 8'h31;
8'h23: output_byte = 8'h32;
8'hc3: output_byte = 8'h33;
8'h18: output_byte = 8'h34;
8'h96: output_byte = 8'h35;
8'h05: output_byte = 8'h36;
8'h9a: output_byte = 8'h37;
8'h07: output_byte = 8'h38;
8'h12: output_byte = 8'h39;
8'h80: output_byte = 8'h3A;
8'he2: output_byte = 8'h3B;
8'heb: output_byte = 8'h3C;
8'h27: output_byte = 8'h3D;
8'hb2: output_byte = 8'h3E;
8'h75: output_byte = 8'h3F;
8'h09: output_byte = 8'h40;
8'h83: output_byte = 8'h41;
8'h2c: output_byte = 8'h42;
8'h1a: output_byte = 8'h43;
8'h1b: output_byte = 8'h44;
8'h6e: output_byte = 8'h45;
8'h5a: output_byte = 8'h46;
8'ha0: output_byte = 8'h47;
8'h52: output_byte = 8'h48;
8'h3b: output_byte = 8'h49;
8'hd6: output_byte = 8'h4A;
8'hb3: output_byte = 8'h4B;
8'h29: output_byte = 8'h4C;
8'he3: output_byte = 8'h4D;
8'h2f: output_byte = 8'h4E;
8'h84: output_byte = 8'h4F;
8'h53: output_byte = 8'h50;
8'hd1: output_byte = 8'h51;
8'h00: output_byte = 8'h52;
8'hed: output_byte = 8'h53;
8'h20: output_byte = 8'h54;
8'hfc: output_byte = 8'h55;
8'hb1: output_byte = 8'h56;
8'h5b: output_byte = 8'h57;
8'h6a: output_byte = 8'h58;
8'hcb: output_byte = 8'h59;
8'hbe: output_byte = 8'h5A;
8'h39: output_byte = 8'h5B;
8'h4a: output_byte = 8'h5C;
8'h4c: output_byte = 8'h5D;
8'h58: output_byte = 8'h5E;
8'hcf: output_byte = 8'h5F;
8'hd0: output_byte = 8'h60;
8'hef: output_byte = 8'h61;
8'haa: output_byte = 8'h62;
8'hfb: output_byte = 8'h63;
8'h43: output_byte = 8'h64;
8'h4d: output_byte = 8'h65;
8'h33: output_byte = 8'h66;
8'h85: output_byte = 8'h67;
8'h45: output_byte = 8'h68;
8'hf9: output_byte = 8'h69;
8'h02: output_byte = 8'h6A;
8'h7f: output_byte = 8'h6B;
8'h50: output_byte = 8'h6C;
8'h3c: output_byte = 8'h6D;
8'h9f: output_byte = 8'h6E;
8'ha8: output_byte = 8'h6F;
8'h51: output_byte = 8'h70;
8'ha3: output_byte = 8'h71;
8'h40: output_byte = 8'h72;
8'h8f: output_byte = 8'h73;
8'h92: output_byte = 8'h74;
8'h9d: output_byte = 8'h75;
8'h38: output_byte = 8'h76;
8'hf5: output_byte = 8'h77;
8'hbc: output_byte = 8'h78;
8'hb6: output_byte = 8'h79;
8'hda: output_byte = 8'h7A;
8'h21: output_byte = 8'h7B;
8'h10: output_byte = 8'h7C;
8'hff: output_byte = 8'h7D;
8'hf3: output_byte = 8'h7E;
8'hd2: output_byte = 8'h7F;
8'hcd: output_byte = 8'h80;
8'h0c: output_byte = 8'h81;
8'h13: output_byte = 8'h82;
8'hec: output_byte = 8'h83;
8'h5f: output_byte = 8'h84;
8'h97: output_byte = 8'h85;
8'h44: output_byte = 8'h86;
8'h17: output_byte = 8'h87;
8'hc4: output_byte = 8'h88;
8'ha7: output_byte = 8'h89;
8'h7e: output_byte = 8'h8A;
8'h3d: output_byte = 8'h8B;
8'h64: output_byte = 8'h8C;
8'h5d: output_byte = 8'h8D;
8'h19: output_byte = 8'h8E;
8'h73: output_byte = 8'h8F;
8'h60: output_byte = 8'h90;
8'h81: output_byte = 8'h91;
8'h4f: output_byte = 8'h92;
8'hdc: output_byte = 8'h93;
8'h22: output_byte = 8'h94;
8'h2a: output_byte = 8'h95;
8'h90: output_byte = 8'h96;
8'h88: output_byte = 8'h97;
8'h46: output_byte = 8'h98;
8'hee: output_byte = 8'h99;
8'hb8: output_byte = 8'h9A;
8'h14: output_byte = 8'h9B;
8'hde: output_byte = 8'h9C;
8'h5e: output_byte = 8'h9D;
8'h0b: output_byte = 8'h9E;
8'hdb: output_byte = 8'h9F;
8'he0: output_byte = 8'hA0;
8'h32: output_byte = 8'hA1;
8'h3a: output_byte = 8'hA2;
8'h0a: output_byte = 8'hA3;
8'h49: output_byte = 8'hA4;
8'h06: output_byte = 8'hA5;
8'h24: output_byte = 8'hA6;
8'h5c: output_byte = 8'hA7;
8'hc2: output_byte = 8'hA8;
8'hd3: output_byte = 8'hA9;
8'hac: output_byte = 8'hAA;
8'h62: output_byte = 8'hAB;
8'h91: output_byte = 8'hAC;
8'h95: output_byte = 8'hAD;
8'he4: output_byte = 8'hAE;
8'h79: output_byte = 8'hAF;
8'he7: output_byte = 8'hB0;
8'hc8: output_byte = 8'hB1;
8'h37: output_byte = 8'hB2;
8'h6d: output_byte = 8'hB3;
8'h8d: output_byte = 8'hB4;
8'hd5: output_byte = 8'hB5;
8'h4e: output_byte = 8'hB6;
8'ha9: output_byte = 8'hB7;
8'h6c: output_byte = 8'hB8;
8'h56: output_byte = 8'hB9;
8'hf4: output_byte = 8'hBA;
8'hea: output_byte = 8'hBB;
8'h65: output_byte = 8'hBC;
8'h7a: output_byte = 8'hBD;
8'hae: output_byte = 8'hBE;
8'h08: output_byte = 8'hBF;
8'hba: output_byte = 8'hC0;
8'h78: output_byte = 8'hC1;
8'h25: output_byte = 8'hC2;
8'h2e: output_byte = 8'hC3;
8'h1c: output_byte = 8'hC4;
8'ha6: output_byte = 8'hC5;
8'hb4: output_byte = 8'hC6;
8'hc6: output_byte = 8'hC7;
8'he8: output_byte = 8'hC8;
8'hdd: output_byte = 8'hC9;
8'h74: output_byte = 8'hCA;
8'h1f: output_byte = 8'hCB;
8'h4b: output_byte = 8'hCC;
8'hbd: output_byte = 8'hCD;
8'h8b: output_byte = 8'hCE;
8'h8a: output_byte = 8'hCF;
8'h70: output_byte = 8'hD0;
8'h3e: output_byte = 8'hD1;
8'hb5: output_byte = 8'hD2;
8'h66: output_byte = 8'hD3;
8'h48: output_byte = 8'hD4;
8'h03: output_byte = 8'hD5;
8'hf6: output_byte = 8'hD6;
8'h0e: output_byte = 8'hD7;
8'h61: output_byte = 8'hD8;
8'h35: output_byte = 8'hD9;
8'h57: output_byte = 8'hDA;
8'hb9: output_byte = 8'hDB;
8'h86: output_byte = 8'hDC;
8'hc1: output_byte = 8'hDD;
8'h1d: output_byte = 8'hDE;
8'h9e: output_byte = 8'hDF;
8'he1: output_byte = 8'hE0;
8'hf8: output_byte = 8'hE1;
8'h98: output_byte = 8'hE2;
8'h11: output_byte = 8'hE3;
8'h69: output_byte = 8'hE4;
8'hd9: output_byte = 8'hE5;
8'h8e: output_byte = 8'hE6;
8'h94: output_byte = 8'hE7;
8'h9b: output_byte = 8'hE8;
8'h1e: output_byte = 8'hE9;
8'h87: output_byte = 8'hEA;
8'he9: output_byte = 8'hEB;
8'hce: output_byte = 8'hEC;
8'h55: output_byte = 8'hED;
8'h28: output_byte = 8'hEE;
8'hdf: output_byte = 8'hEF;
8'h8c: output_byte = 8'hF0;
8'ha1: output_byte = 8'hF1;
8'h89: output_byte = 8'hF2;
8'h0d: output_byte = 8'hF3;
8'hbf: output_byte = 8'hF4;
8'he6: output_byte = 8'hF5;
8'h42: output_byte = 8'hF6;
8'h68: output_byte = 8'hF7;
8'h41: output_byte = 8'hF8;
8'h99: output_byte = 8'hF9;
8'h2d: output_byte = 8'hFA;
8'h0f: output_byte = 8'hFB;
8'hb0: output_byte = 8'hFC;
8'h54: output_byte = 8'hFD;
8'hbb: output_byte = 8'hFE;
8'h16: output_byte = 8'hFF;
endcase
end
endmodule